module main

import mymodule

fn main() {
    mymodule.say_hi()
}
