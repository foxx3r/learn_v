module mymodule

pub fn say_hi() {
    println("Hello from mymodule!")
}
